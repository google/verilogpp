// busthing

module busthing #(
  parameter WIDTH = 5
) (
  input logic [WIDTH-1:0] i
);

foo i foo

endmodule

