module drive_two (
  output logic [1:0] foo
);

assign foo = 1'b1;

endmodule : drive_one
