module drive_one(
  output logic foo
);

assign foo = 1'b1;

endmodule : drive_one
